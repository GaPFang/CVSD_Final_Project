`include "../01_RTL/ed25519.sv"
`include "../01_RTL/scalarMul_wNAF_Extended.sv"
`include "../01_RTL/pointAddExtended.sv"
`include "../01_RTL/numberMul.sv"
`include "../01_RTL/reduction.sv"
`include "../01_RTL/montgomeryInv.sv"
